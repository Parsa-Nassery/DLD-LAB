library verilog;
use verilog.vl_types.all;
entity transTB is
end transTB;
