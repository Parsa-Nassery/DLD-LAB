module Adder(input [7:0] a, input b, output [7:0]out);
	assign out = a + b + 1;
endmodule