library verilog;
use verilog.vl_types.all;
entity SSDTB is
end SSDTB;
