library verilog;
use verilog.vl_types.all;
entity TBOnePulser is
end TBOnePulser;
