library verilog;
use verilog.vl_types.all;
entity EXPTB is
end EXPTB;
